//--------------------------------------------------------------------
// Design Name : core
// File Name   : core.sv
// Function    :  
// Designer    : Chen Xiaowei         - Nanyang technological University 
//                                    - Technische Universität München
// Email       : chen1408@e.ntu.edu.sg
// Blog         : haitianzhishang.github.io
//---------------------------------------------------------------------
module core #(
  parameter  
)
(
  input             clk,    
  input             rst_n, 
  input    [  :  ]    ,
  output   [  :  ]    ,
  
);

always@(posedge clk or negedge rst) 
begin
  if(!rst) 
  begin
    
  end
  else
  begin
    
  end
end

always@(*) 
begin

end

endmodule : core